library verilog;
use verilog.vl_types.all;
entity ControlAscensor_vlg_vec_tst is
end ControlAscensor_vlg_vec_tst;
