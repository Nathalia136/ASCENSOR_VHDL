library verilog;
use verilog.vl_types.all;
entity ContadorPersonas_vlg_vec_tst is
end ContadorPersonas_vlg_vec_tst;
