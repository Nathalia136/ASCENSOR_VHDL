library verilog;
use verilog.vl_types.all;
entity ControladorPuertas_vlg_vec_tst is
end ControladorPuertas_vlg_vec_tst;
