library verilog;
use verilog.vl_types.all;
entity gestion_cabina_vlg_vec_tst is
end gestion_cabina_vlg_vec_tst;
