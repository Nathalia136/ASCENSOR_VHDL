library verilog;
use verilog.vl_types.all;
entity identificador_direccion_vlg_vec_tst is
end identificador_direccion_vlg_vec_tst;
