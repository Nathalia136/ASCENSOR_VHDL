library verilog;
use verilog.vl_types.all;
entity gestion_externas_vlg_vec_tst is
end gestion_externas_vlg_vec_tst;
