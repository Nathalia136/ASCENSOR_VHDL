library verilog;
use verilog.vl_types.all;
entity ControladorPuertas_vlg_check_tst is
    port(
        puerta          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ControladorPuertas_vlg_check_tst;
