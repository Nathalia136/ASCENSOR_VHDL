library verilog;
use verilog.vl_types.all;
entity Alarmas_vlg_vec_tst is
end Alarmas_vlg_vec_tst;
