library verilog;
use verilog.vl_types.all;
entity detectar_piso_actual_vlg_vec_tst is
end detectar_piso_actual_vlg_vec_tst;
